package profiler_dpi_pkg;
  `include "profiler_dpi.svh"
endpackage
