`ifndef INCLUDED_srm_base_observer
`define INCLUDED_srm_base_observer

virtual class srm_base_observer;
  pure virtual function void sample(const ref srm_generic_xact_t xact); 
endclass

`endif
