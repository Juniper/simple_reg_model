// Package for unit test framework
`ifndef INCLUDED_srm_unit_test_pkg
`define INCLUDED_srm_unit_test_pkg

package srm_unit_test_pkg;
  `include "srm_unit_test.svh"
endpackage

`endif
